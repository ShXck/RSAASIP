module sum(input logic[28:0] a, b, output logic[28:0] out);

assign out = a + b;

endmodule
